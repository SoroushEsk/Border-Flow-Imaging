`timescale 1ns / 1ps



module FPGA_Sender(
							input clk
    );


endmodule
