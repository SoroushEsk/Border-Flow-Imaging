`timescale 1ns / 1ps

`define Initial 0
`define StartPoint 1
`define FindCode 2
`define FindArea 3
`define DoneAnalysing 4

module FPGA_Reciever(
	input clk
    );


endmodule
