module FPGA_Reciever(
	input clk
    );


endmodule
