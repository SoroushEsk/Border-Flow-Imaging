`timescale 1ns / 1ps



module FPGA_Sender(
							input Clk, 
							input reset,
							output UART_Out
    );


endmodule
